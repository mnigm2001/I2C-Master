`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/07/2025 10:04:29 PM
// Design Name: 
// Module Name: i2c_master_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module i2c_master_tb();

//    clk_divider_tb clk_divider_test();

/*
input wire clk,
    input wire resetn,
    input wire start,
    output reg busy,
    output reg [15:0] data_out,
    output reg data_valid,
    inout wire sda

input wire clk,
    input wire resetn,
    input wire start,
    output reg busy,
    output reg [15:0] data_out,
    output reg data_valid,
    output reg scl,
    inout wire sda
    
*/

    
    localparam SLAVE_ADDR = 7'b1001000;
    
    /* Master Ports */
    logic clk=0;
    logic resetn;
    
    logic start;
    logic busy;
    logic [15:0] data_out;
    logic data_valid;
    wire sda;  // inout
    logic scl;
    
    i2c_master DUT (
        .clk(clk),
        .resetn(resetn),
        .start(start),
        .busy(busy),
        .data_out(data_out),
        .data_valid(data_valid),
        .scl(scl),
        .sda(sda)
    );
    
    /* Slave Ports */
    logic clk_sl=0;
//    logic scl;
    
    // Generate master CLK
    always #10 clk = ~clk;
    
    // Generate slave CLK (for simulation purposes) -- actual clock actually generated by master
    always #5000 clk_sl = ~clk_sl;
    
    /*
        50Mhz at 1ns/1ps
        frequency = nEm
        delay = ((1/nEm)/timescale)/2
        
        100khz at 1ns
        delay = 5000
    
    */
    
    initial begin
    
        start = 1'b0;
    
        resetn = 1'b1;
        @(posedge clk);
        resetn = 1'b0;
        repeat (3) @(posedge clk);
        resetn = 1'b1;
        #500;
        
        // Start
        @(posedge clk);
        start = 1'b1;
        
        // Addr
        @(posedge clk);
        start = 1'b0;
        repeat (10) @(posedge clk_sl);

        
        
        
        
        #1000;
        $finish;
    end
    
    
    
    
    
    

    
//    task master_write(input [6:0] addr, input [7:0] data, inout sda, output scl);
//        if (start) begin
//            sda = 1'b0; // Start
//            scl = 1'b0;
//        end
//        // 
//        for (int i=0; i<8; i++) begin
//            repeat (250) @(posedge clk);
//            scl = 1'b1; 
            
//        end
////    send_byte({addr, 1'b0});
////    wait_for_ack();
////    send_byte(data);
////    wait_for_ack();
////    send_stop();


//    endtask
    
    
////    task slave_read(input scl, inout sda);
        
////    endtask
endmodule






//    task gen_scl(input en, output scl);
//        scl = 1'b1;
//        if (en) begin
//            #10 scl = ~scl; 
//        end
//    endtask




